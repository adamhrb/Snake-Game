
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; -- Use numeric_std instead of std_logic_unsigned

entity Basic_ROM is
    Port ( addr : in  STD_LOGIC_VECTOR (4 downto 0);
           M : out  STD_LOGIC_VECTOR (11 downto 0));
end Basic_ROM;

architecture Behavioral of Basic_ROM is
type rom_array is array (NATURAL range <>) of std_logic_vector(11 downto 0);

--constant rom:rom_array:= (
--	"111111111111", "111111111111", "111111111111", "111111111111","111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", --0 --> 15
--	"111111111111", "111111111111", "111111111111", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "111111111111", "111111111111", "111111111111", --16 --> 31
--	"111111111111", "111111111111", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "111111111111", --32 --> 47
--	"111111111111", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000","000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", --48 --> 63
--	"111111111111", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000","000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "111111111111", --64 --> 79
--	"000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", --80 --> 95
--	"000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", --96 --> 111
--	"000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", --112 --> 127
--	"000000000000", "000000000000", "000000000000", "000000000000","000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111","111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", --128 --> 139
--	"000000000000", "000000000000", "000000000000", "000000000000","000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111","111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", --140 --> 159 
--	"000000000000", "000000000000", "000000000000", "000000000000","111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111","111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", --160 --> 175
--	"111111111111", "000000000000", "000000000000", "000000000000","111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000","111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "111111111111", --176 --> 191
--	"111111111111", "000000000000", "000000000000", "000000000000","111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000","111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "111111111111", --192 --> 207
--	"111111111111", "111111111111", "000000000000", "000000000000","000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111","111111111111", "111111111111", "000000000000", "000000000000", "111111111111", "111111111111", --208 --> 223
--	"111111111111", "111111111111", "111111111111", "000000000000","000000000000", "000000000000", "000000000000", "111111111111", "111111111111", "111111111111","111111111111", "000000000000", "000000000000", "111111111111", "111111111111", "111111111111", --224 --> 239
--	"111111111111", "111111111111", "111111111111", "111111111111","111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000","000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"  --240 --> 255 
--	);

constant rom:rom_array:= (
	"111111111111", "111111111111", "111111111111", "111111111111", --0 --> 3
	"111111111111", "000000000000", "000000000000", "111111111111", --4 --> 7
	"111111111111", "000000000000", "000000000000", "111111111111", --8 --> 11
	"111111111111", "000000000000", "000000000000", "111111111111", --12 --> 15
	"111111111111", "111111111111", "111111111111", "111111111111" --16 --> 19
	);
	
begin

process(addr)
variable j: integer;

begin
	j := to_integer(unsigned(addr)); -- Convert using numeric_std
	if (j < 20) then M <= rom(j);
	else M <= (others =>'0');
	end if;

end process;
end Behavioral;
